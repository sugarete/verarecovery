module XTS (
    input [0:127] key1,
    input [0:127] key2,
    input [0:127] data,
    input [0:127] tweak,
    output [0:127] result
);

//---------wires, registers----------    


endmodule