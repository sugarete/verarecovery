module Decrypt_Serpent (
    input wire [255:0] i_key,
    input wire [127:0] i_data,
    output wire [127:0] o_data
);
    
endmodule